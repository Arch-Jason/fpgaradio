// cordic.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module cordic (
		input  wire [11:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [7:0]  c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [7:0]  s       //      s.s
	);

	cordic_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
